
  //------------------------------------//
 //            TIME                    //
//------------------------------------//
/*------------------------------------------------------------------------------                    
    freq
-------------------------------------------------------------------------------*/ 
localparam   SYS_CLK_FREQ = 74 ; //*100kHz

localparam   TIME_0P5uS  = SYS_CLK_FREQ / 20       ;
localparam   TIME_1uS    = SYS_CLK_FREQ / 10       ;
localparam   TIME_2uS    = SYS_CLK_FREQ / 5        ;
localparam   TIME_3uS    = SYS_CLK_FREQ / 3        ;
localparam   TIME_5uS    = SYS_CLK_FREQ / 2        ;
localparam   TIME_10uS   = SYS_CLK_FREQ            ;
localparam   TIME_20uS   = SYS_CLK_FREQ * 2        ;
localparam   TIME_50uS   = SYS_CLK_FREQ * 5        ;
localparam   TIME_100uS  = SYS_CLK_FREQ * 10       ;
localparam   TIME_150uS  = SYS_CLK_FREQ * 15       ;

localparam   TIME_1mS    = SYS_CLK_FREQ * 100      ;
localparam   TIME_5mS    = SYS_CLK_FREQ * 500      ;
localparam   TIME_10mS   = SYS_CLK_FREQ * 1000     ;
localparam   TIME_300mS  = SYS_CLK_FREQ * 30000    ;
localparam   TIME_400mS  = SYS_CLK_FREQ * 40000    ;

localparam   TIME_2S     = SYS_CLK_FREQ * 200000   ;





