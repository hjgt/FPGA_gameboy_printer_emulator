function integer clogb2 (input integer size);
  begin
    size = size - 1;
    for (clogb2=1; size>1; clogb2=clogb2+1)
      size = size >> 1;
  end
endfunction // clogb2